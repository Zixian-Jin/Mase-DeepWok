/*
 * fixed_linear_sparse: matmul(data_in, weight)
 * Three trucks in each row of weight are streamed together at every clock cycle
 * Assumption: two trucks out of tree are always sparse
 * Expected throughput: every IN_DEPTH/3 cycles. i.e., 3x speed up compared with fixed_linear.sv 
 */
`timescale 1ns / 1ps
module fixed_linear_sparse #(
    /* sparsity-related params */
    parameter BLOCK_SIZE = 4,
    parameter WEIGHT_BLOCKS = 3,
    parameter WEIGHT_BLOCKS_SPARSE = 2,

    parameter IN_WIDTH = 32,
    parameter IN_FRAC_WIDTH = 0,
    parameter IN_SIZE = BLOCK_SIZE * WEIGHT_BLOCKS,
    parameter IN_DEPTH = 3,
    parameter PARALLELISM = 2,

    parameter WEIGHT_WIDTH = 16,
    parameter WEIGHT_FRAC_WIDTH = 0,
    parameter WEIGHT_SIZE = BLOCK_SIZE * WEIGHT_BLOCKS * PARALLELISM,


    // This is the width for the summed product
    // +1 is because of the bias
    parameter HAS_BIAS = 0,
    parameter OUT_WIDTH = IN_WIDTH + WEIGHT_WIDTH + $clog2(BLOCK_SIZE*(WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE)) + $clog2(IN_DEPTH) + HAS_BIAS,
    /* verilator lint_off UNUSEDPARAM */
    parameter OUT_FRAC_WIDTH = IN_FRAC_WIDTH + WEIGHT_FRAC_WIDTH,
    /* verilator lint_on UNUSEDPARAM */
    parameter OUT_SIZE = PARALLELISM,

    parameter BIAS_SIZE = OUT_SIZE,
    parameter BIAS_WIDTH = 32,
    /* verilator lint_off UNUSEDPARAM */
    parameter BIAS_FRAC_WIDTH = 0
    /* verilator lint_on UNUSEDPARAM */
) (
    input clk,
    input rst,

    // input port for data_inivations
    input  [IN_WIDTH-1:0] data_in      [IN_SIZE-1:0],
    input                 data_in_valid,
    output                data_in_ready,

    // input port for weight
    input  [WEIGHT_WIDTH-1:0] weight      [WEIGHT_SIZE-1:0],
    input                     weight_valid,
    output                    weight_ready,

    /* verilator lint_off UNUSEDSIGNAL */
    input  [BIAS_WIDTH-1:0] bias          [BIAS_SIZE-1:0],
    input                   bias_valid,
    /* verilator lint_on UNUSEDSIGNAL */
    output                  bias_ready,
    output [ OUT_WIDTH-1:0] data_out      [ OUT_SIZE-1:0],
    output                  data_out_valid,
    input                   data_out_ready
);

  localparam FDP_WIDTH = IN_WIDTH + WEIGHT_WIDTH + $clog2(BLOCK_SIZE*(WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE));
  localparam ACC_WIDTH = FDP_WIDTH + $clog2(IN_DEPTH);

  logic fdp_join_valid, fdp_join_ready;
  join2 #() fdp_join_inst (
      .data_in_ready ({weight_ready, data_in_ready}),
      .data_in_valid ({weight_valid, data_in_valid}),
      .data_out_valid(fdp_join_valid),
      .data_out_ready(fdp_join_ready)
  );

  /* verilator lint_off UNUSEDSIGNAL */
  // Assume the parallelised hardware above have the same arrival time
  // which means that they always have the same state. So we can just
  // pick one of the valid signal to use.
  logic [PARALLELISM-1:0] fdp_data_ready, fdp_weight_ready;
  assign fdp_join_ready = fdp_data_ready[0];
  /* verilator lint_on UNUSEDSIGNAL */

  logic                 acc_ready;
  logic [ACC_WIDTH-1:0] acc_data_out[PARALLELISM-1:0];




  // There are PARALLELISM number of dot product instances with IN_SIZE inputs 
  // and each one computes for IN_DEPTH iterations for each inputs.
  for (genvar i = 0; i < PARALLELISM; i = i + 1) begin : linear
    // Assume the weight are transposed and partitioned 
    logic [WEIGHT_WIDTH-1:0] current_weight[IN_SIZE-1:0];
    assign current_weight = weight[IN_SIZE*(i+1)-1:IN_SIZE*i];

    /* sparsity related logics */
    logic [WEIGHT_BLOCKS-1:0] nzc_result;
    logic [WEIGHT_WIDTH-1:0] current_active_weight[BLOCK_SIZE*(WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE)-1 : 0];
    logic [IN_WIDTH-1:0] current_active_data_in[BLOCK_SIZE*(WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE)-1 : 0];
    // localparam NON_ZERO_INDEX = 0; // assume only the first block is non-sparse
    // logic [31:0] non_zero_block_id;
    // logic [31:0] non_zero_blocks;  // assumed to be constant

    for (genvar j = 0; j < WEIGHT_BLOCKS; j = j + 1) begin: NZC
        nzc #(
            .IN_WIDTH (WEIGHT_WIDTH),
            .IN_SIZE (BLOCK_SIZE)
        ) nzc_inst (
            .data_in (current_weight[BLOCK_SIZE*(j+1)-1: BLOCK_SIZE*j]),
            .zero_flag (nzc_result[j])
        );

        // always_comb begin
        //     /* verilator lint_off LATCH */
        //     if (zero_flag) begin
        //         current_active_weight = current_weight[BLOCK_SIZE*(j+1)-1: BLOCK_SIZE*j];
        //         current_active_data_in = data_in[BLOCK_SIZE*(j+1)-1: BLOCK_SIZE*j];
        //     end
            // else begin
            //     current_active_weight = current_active_weight;
            //     current_active_data_in = current_active_data_in;
            // end
        // end
    end

    MUX #(
        .IN_BLOCK_NUM (WEIGHT_BLOCKS),
        .BLOCK_SIZE (BLOCK_SIZE),
        .OUT_BLOCK_NUM (WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE),
        .IN_WIDTH (WEIGHT_WIDTH)
    ) mux_inst_weight (
        .nonzero_sel (nzc_result),
        .din (current_weight),
        .dout (current_active_weight)
    );

    MUX #(
        .IN_BLOCK_NUM (WEIGHT_BLOCKS),
        .BLOCK_SIZE (BLOCK_SIZE),
        .OUT_BLOCK_NUM (WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE),
        .IN_WIDTH (IN_WIDTH)
    ) mux_inst_data_in (
        .nonzero_sel (nzc_result),
        .din (data_in),
        .dout (current_active_data_in)
    );
    // for (genvar k = 0; k < WEIGHT_BLOCKS; k = k + 1) begin
    //     always_comb begin
    //         if (nzc_result[k] == 1'b0) begin
    //             current_active_weight = current_weight[BLOCK_SIZE*(k+1)-1: BLOCK_SIZE*k];
    //             current_active_data_in = data_in[BLOCK_SIZE*(k+1)-1: BLOCK_SIZE*k];
    //         end
    //         else begin
    //             current_active_weight = current_weight[BLOCK_SIZE*(k+1)-1: BLOCK_SIZE*k];
    //             current_active_data_in = data_in[BLOCK_SIZE*(k+1)-1: BLOCK_SIZE*k];
    //         end
    //     end
    // end
    // assign current_active_weight = current_weight[BLOCK_SIZE*(NON_ZERO_INDEX+1)-1: BLOCK_SIZE*NON_ZERO_INDEX];
    // assign current_active_data_in = data_in[BLOCK_SIZE*(NON_ZERO_INDEX+1)-1: BLOCK_SIZE*NON_ZERO_INDEX];

    logic [FDP_WIDTH-1:0] fdp_data_out;
    logic fdp_data_out_valid, fdp_data_out_ready;

    // The inputs are already sync-ed by the previous join
    fixed_dot_product #(
        .IN_WIDTH(IN_WIDTH),
        .WEIGHT_WIDTH(WEIGHT_WIDTH),
        .IN_SIZE(BLOCK_SIZE*(WEIGHT_BLOCKS-WEIGHT_BLOCKS_SPARSE))
    ) fdp_inst (
        .clk(clk),
        .rst(rst),
        .data_in(current_active_data_in),
        .data_in_valid(fdp_join_valid),
        .data_in_ready(fdp_data_ready[i]),
        .weight(current_active_weight),
        .weight_valid(fdp_join_valid),
        .weight_ready(fdp_weight_ready[i]),
        .data_out(fdp_data_out),
        .data_out_valid(fdp_data_out_valid),
        .data_out_ready(fdp_data_out_ready)
    );

    /* verilator lint_off UNUSEDSIGNAL */
    logic acc_data_out_valid, acc_data_out_ready;
    /* verilator lint_on UNUSEDSIGNAL */


    // /* NZC-gating for sparse vector computation */
    logic zero_flag;
    assign zero_flag = 1'b0;
    logic [FDP_WIDTH-1:0] acc_data_in;
    logic acc_data_in_valid, acc_data_in_ready;

    // always_comb begin
    //     if (data_in[0] == 0 || data_in[1] == 0 || data_in[2] == 0 || data_in[3] == 0) zero_flag = 1'b1;
    //     else if (current_weight[0] == 0 || current_weight[1] == 0 || current_weight[2] == 0 || current_weight[3] == 0) zero_flag = 1'b1;
    //     else zero_flag = 1'b0;
    // end

    assign acc_data_in = zero_flag ? 0 : fdp_data_out;
    assign acc_data_in_valid = zero_flag ? 1 : fdp_data_out_valid;
    assign fdp_data_out_ready = zero_flag ? 0 : acc_data_in_ready; 

    fixed_accumulator #(
        .IN_WIDTH(FDP_WIDTH),
        .IN_DEPTH(IN_DEPTH)
    ) fixed_accumulator_inst (
        .clk(clk),
        .rst(rst),
        .data_in(acc_data_in),
        .data_in_valid(acc_data_in_valid),
        .data_in_ready(acc_data_in_ready),
        .data_out(acc_data_out[i]),
        .data_out_valid(acc_data_out_valid),
        .data_out_ready(acc_data_out_ready)
    );

    // Assume the parallelised hardware above have the same arrival time
    // which means that they always have the same state. So we can just
    // pick one of the valid signal to use.
    assign acc_data_out_ready = acc_ready;
  end


  if (HAS_BIAS == 1) begin

    logic [ACC_WIDTH-1:0] bias_sext[PARALLELISM-1:0];
    join2 #() acc_join_inst (
        .data_in_ready ({bias_ready, acc_ready}),
        .data_in_valid ({bias_valid, linear[0].acc_data_out_valid}),
        .data_out_valid(acc_join_valid),
        .data_out_ready(acc_join_ready)
    );
    logic [PARALLELISM-1:0] reg_ready;
    assign acc_join_ready = &reg_ready;

    logic acc_join_valid, acc_join_ready;
    fixed_rounding #(
        .IN_SIZE(PARALLELISM),
        .IN_WIDTH(BIAS_WIDTH),
        .IN_FRAC_WIDTH(BIAS_FRAC_WIDTH),
        .OUT_WIDTH(ACC_WIDTH),
        .OUT_FRAC_WIDTH(IN_FRAC_WIDTH + WEIGHT_FRAC_WIDTH)
    ) bias_cast (
        .data_in (bias),
        .data_out(bias_sext)
    );

    for (genvar i = 0; i < PARALLELISM; i = i + 1) begin : add_bias
      logic [OUT_WIDTH-1:0] add;
      assign add = $signed(acc_data_out[i]) + $signed(bias_sext[i]);
      /* verilator lint_off UNUSEDSIGNAL */
      logic dout_valid;
      skid_buffer #(
          .DATA_WIDTH(OUT_WIDTH)
      ) register_slice (
          .clk           (clk),
          .rst           (rst),
          .data_in_valid (acc_join_valid),
          .data_in_ready (reg_ready[i]),
          .data_in       (add),
          .data_out_valid(dout_valid),
          .data_out_ready(data_out_ready),
          .data_out      (data_out[i])
      );
    end
    assign data_out_valid = add_bias[0].dout_valid;

  end else begin
    assign acc_ready = data_out_ready;
    assign data_out_valid = linear[0].acc_data_out_valid;
    assign data_out = acc_data_out;
    assign bias_ready = 1;
  end

endmodule
